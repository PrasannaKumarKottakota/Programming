`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 5G Testbed, IISc
// Engineer: K. Prasanna Kumar 
// Module Name: SR_LATCH_tb
//////////////////////////////////////////////////////////////////////////////////


module SR_LATCH_tb(

    );
endmodule
