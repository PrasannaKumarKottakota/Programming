`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 5G Testbed, IISc 
// Engineer: K. Prasanna Kumar
// Module Name: D_flipflop
//////////////////////////////////////////////////////////////////////////////////


module D_flipflop(D, Q, Q_bar);
input D;
output Q, Q_bar;

sr_latch SRL (D, ~D, Q, Q_bar);

endmodule
