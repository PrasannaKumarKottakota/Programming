`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: IISc 
// Engineer: K. Prasanna Kumar
// 
//////////////////////////////////////////////////////////////////////////////////


module sr_latch(R, S, Q, Qbar);
input R, S;
output Q, Qbar;

assign Q = ~(R & Qbar);
assign Qbar = ~(S & Q);
endmodule
